`include  "memoria.v"

module bancoPrueba;



true_dpram_sclk memoria (
    //OUTPUTS
    .q_a    (),
    .q_b    (),
    //INPUTS
    .data_a (),
    .data_b (),
    .addr_a (),
    .addr_b (),
    .we_a   (),
    .we_b   (),
    .clk    ()
);

probador probador1(







);


endmodule